// Generator : SpinalHDL v1.6.2    git head : 6f25d9a541c42028018402843d80c1b0948f0d13
// Component : Wire_1

`timescale 1ns/1ps 

module Wire_1 (
  input      [0:0]    io_i,
  output     [0:0]    io_o
);


  assign io_o = io_i;

endmodule
